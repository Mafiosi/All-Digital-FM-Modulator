/*
    Spartan 6 board testbench for PSD2018/2019 lab3 project (V1.0 - 26 Dec 2018)
	
    jca@fe.up.pt

	This Verilog code is property of University of Porto
	Its utilization beyond the scope of the course Digital Systems Design
	(Projeto de Sistemas Digitais) of the Integrated Master in Electrical 
	and Computer Engineering requires explicit authorization from the author.
	
*/
`timescale 1ns/1ps

// Configure testbench: Uncomment the following 'define' to enable debugging:
`define DEBUG_PRINT         // Print NDATA_TO_PRINT correct or error results
`define NDATA_TO_PRINT 20   // Number of OK/NOK results to print

/* KEEP THIS HERE BUT DO NOT USE IN THIS TESTBENCH
// `define DEBUG_PROBES   5   // Print the first N results at each 192k and 48k clock cycles:
*/

// Number of input samples to simulate
// set this constant to a constant integer or to the variable 'no_input_samples' that
// will be loaded with the actual number of input samples read from the input audio files
`define NSAMPLES_SIM   no_input_samples


module s6base_tb;

//--------------------------------------------------------------------
// primary inputs:								
// clocks:
reg				clk100M, reset_n;

// push buttons:
wire				btnu, btnr, btnd, btnl, btnc;
reg       [4:0]     btns;

// slide switches:
wire				sw7, sw6, sw5, sw4, sw3, sw2, sw1, sw0;
reg       [7:0]     sws;

// LEDs:
wire 			    ld0, ld1, ld2, ld3, ld4, ld5, ld6, ld7;
wire      [7:0]     leds;

// RS232:
wire			rx, tx;

// LM4450 audio CODEC:
// These signals are driven by the LM4550 verification IP
reg  XTAL_IN;
wire RESET_N, SYNC;
wire SDATA_OUT;
wire BIT_CLK, SDATA_IN;

// PMOD connector (to the DAC):
wire PMOD1, PMOD2, PMOD3, PMOD4, PMOD7, PMOD8, PMOD9, PMOD10;


// VHDC connector:
wire VHDC1P,  VHDC1N, VHDC2P, VHDC2N, VHDC3P, VHDC3N, VHDC4P, VHDC4N, 
     VHDC5P,  VHDC5N, VHDC6P, VHDC6N, VHDC7P, VHDC7N, VHDC8P, VHDC8N, 
     VHDC9P,  VHDC9N,  VHDC10P, VHDC10N, VHDC11P, VHDC11N, VHDC12P, VHDC12N,
     VHDC13P, VHDC13N, VHDC14P, VHDC14N, VHDC15P, VHDC15N, VHDC16P, VHDC16N,
     VHDC17P, VHDC17N, VHDC18P, VHDC18N, VHDC19P, VHDC19N, VHDC20P, VHDC20N;


	 
// -----------------------------------------------------------------
// Testbench configuration parameters:         
parameter           
          // audio input files created by the Matlab script 'fmstereo_gensimdata.m'
          LEFT_IN_FILENAME  = "../simdata/fmstereo_audioin_left.hex",
		  RIGHT_IN_FILENAME = "../simdata/fmstereo_audioin_right.hex",
		  
		  // The file generated by the same script with the golden results
		  // at the output of the FM stereo encoder, before the final DDS:
		  FM_GOLDEN_OUTPUT_FILENAME  = "../simdata/fmstereo_mpx_golden.hex",
		  DAC_GOLDEN_OUTPUT_FILENAME = "../simdata/DAC_golden.hex",

          // The output files created by the simulation. 
		  FM_OUTPUT_FILENAME    = "../simdata/fmstereo_mpx.hex",
		  DAC_OUTPUT_FILENAME   = "../simdata/DACoutput.hex",

		  // Input parameters:
          FREQ_STEPWC = 18'b000010001001010100, // stepWC, FM freqs 95.50 ans 101.60 MHz
		  GAIN_Ks = 4'b0_100,     //     0.100b = 0.5 decimal
          GAIN_Kd = 4'b1_000,     //     1.000b = 1.0 decimal
          GAIN_Kp = 4'b0_001,     //     0.100b = 0.5 decimal
          GAIN_Kf = 8'b0100_0000, // 0100.0000b = 4.0 decimal
		  
		  MAX_ERRORS          = 20,             // Number of errors found that will stop the simulation
		  
		  // Set the maximum simulation time, as the number of input sampling periods
		  // or approximately number of input samples. 
		  // Simulation stops when this time is exhausted or when input samples end
		  MAX_SIMULATION_TIME = 48_000*1,       // This simulates only 1 second of real time	

//###########################################################################################################
// DO NOT TOUCH BELOW THIS LINE ** DO NOT TOUCH BELOW THIS LINE ** DO NOT TOUCH BELOW THIS LINE ** 		  
//###########################################################################################################
		  
		  CLOCKS_PER_SAMPLE  = 256,              // Number of clock cycles per input sampling period
		  MAX_INPUT_SIZE     = 48000 * 2,        // max number of samples of input audio files (2 == 2 seconds)

          // Configure testbench clocks: The design is driven by BIT_CLK (12.288 MHz) generated by
		  // the audio codec. This signal is derived from a 24.576 MHz oscillator 
		  CLOCK_FREQUENCY    = 48000 * CLOCKS_PER_SAMPLE,     // Bit clock, Hertz (12.288 MHz)
		  CLOCK_PERIOD       = 1/CLOCK_FREQUENCY,             // seconds
		  CLOCK_PERIOD_NS    = 1000000000.0/CLOCK_FREQUENCY,    // clock period, in nanoseconds
		  
		  // The external oscillator:
		  XTAL_FREQUENCY     = 48000 * CLOCKS_PER_SAMPLE * 2, // 24.576 MHz
		  XTAL_PERIOD_NS     = 1000000000.0/XTAL_FREQUENCY,   //clock period in ns
		  
		  INTERNAL_CLOCK_PERIOD = 1000000000.0/( CLOCK_FREQUENCY * 8.0 ), // Internal master clock
		  
		  N_SAMPLES_LATENCY     = 3, // Latency of the audio CODEC simulation model (# of sampling periods)
		  
 		  N_CLOCKS_RESET  = 2;                  // Number of clock cycles for applying reset



s6base s6base_1( 
				//------------------------------------------------------------------
                // external clock source:
               .clockext100MHz(clk100M),	// master clock input (external oscillator 100MHz)
               .reset_n(reset_n),           // external reset, active low
				//------------------------------------------------------------------
                // push buttons: button down = logic 1 (no debouncing hw)
				.btnu( btnu ),			// button up
				.btnr( btnr ),
				.btnd( btnd ),
				.btnl( btnl ),			// button left
				.btnc( btnc ),          // button center

				//------------------------------------------------------------------
                // Slide switches:
				.sw0( sw0 ),
				.sw1( sw1 ),
				.sw2( sw2 ),
				.sw3( sw3 ),
				.sw4( sw4 ),
				.sw5( sw5 ),
				.sw6( sw6 ),
				.sw7( sw7 ),

				//------------------------------------------------------------------
				// LEDs: logic 1 lights the LED
				.ld7( ld7 ),			// LED 7 (leftmost)
				.ld6( ld6 ),
				.ld5( ld5 ),
				.ld4( ld4 ),
				.ld3( ld3 ),
				.ld2( ld2 ),
				.ld1( ld1 ),
				.ld0( ld0 ),			// LED 0 (rightmost)


				//------------------------------------------------------------------
				// Serial interface (RS232 port)
               .tx( tx ),			// tx data (output from the user circuit)
               .rx( rx ),
				
				//------------------------------------------------------------------	 
				// Audio codec interface (AC97)
				.SDATA_IN(SDATA_IN),
				.SDATA_OUT(SDATA_OUT),
				.SYNC(SYNC),
				.BIT_CLK(BIT_CLK),
				.RESET_N(RESET_N),
				
			    //------------------------------------------------------------------
			    // PMOD connector
			   .PMOD1(  PMOD1 ),  
			   .PMOD2(  PMOD2 ),  
			   .PMOD3(  PMOD3 ),  
			   .PMOD4(  PMOD4 ),  
			   .PMOD7(  PMOD7 ),  
			   .PMOD8(  PMOD8 ),  
			   .PMOD9(  PMOD9 ),  
			   .PMOD10( PMOD10 ),
			   
			   // VHDC connector
			   .VHDC1P(  VHDC1P ),
			   .VHDC1N(  VHDC1N ),
			   .VHDC2P(  VHDC2P ),
			   .VHDC2N(  VHDC2N ),
			   .VHDC3P(  VHDC3P ),
			   .VHDC3N(  VHDC3N ),
			   .VHDC4P(  VHDC4P ),
			   .VHDC4N(  VHDC4N ),
			   .VHDC5P(  VHDC5P ),
			   .VHDC5N(  VHDC5N ),
			   .VHDC6P(  VHDC6P ),
			   .VHDC6N(  VHDC6N ),
			   .VHDC7P(  VHDC7P ),
			   .VHDC7N(  VHDC7N ),
			   .VHDC8P(  VHDC8P ),
			   .VHDC8N(  VHDC8N ),
			   .VHDC9P(  VHDC9P ),
			   .VHDC9N(  VHDC9N ),
			   .VHDC10P( VHDC10P ),
			   .VHDC10N( VHDC10N ),
			   .VHDC11P( VHDC11P ),
			   .VHDC11N( VHDC11N ),
			   .VHDC12P( VHDC12P ),
			   .VHDC12N( VHDC12N ),
			   .VHDC13P( VHDC13P ),
			   .VHDC13N( VHDC13N ),
			   .VHDC14P( VHDC14P ),
			   .VHDC14N( VHDC14N ),
			   .VHDC15P( VHDC15P ),
			   .VHDC15N( VHDC15N ),
			   .VHDC16P( VHDC16P ),
			   .VHDC16N( VHDC16N ),
			   .VHDC17P( VHDC17P ),
			   .VHDC17N( VHDC17N ),
			   .VHDC18P( VHDC18P ),
			   .VHDC18N( VHDC18N ),
			   .VHDC19P( VHDC19P ),
			   .VHDC19N( VHDC19N ),
			   .VHDC20P( VHDC20P ),
			   .VHDC20N( VHDC20N )         			 
);

// VHDC bus (for routing signals to primary outputs):
// assign unused outputs to zero.
wire [39:0] VHDC = 
   { VHDC1P,  VHDC1N, VHDC2P, VHDC2N, VHDC3P, VHDC3N, VHDC4P, VHDC4N, 
     VHDC5P,  VHDC5N, VHDC6P, VHDC6N, VHDC7P, VHDC7N, VHDC8P, VHDC8N, 
     VHDC9P,  VHDC9N,  VHDC10P, VHDC10N, VHDC11P, VHDC11N, VHDC12P, VHDC12N,
     VHDC13P, VHDC13N, VHDC14P, VHDC14N, VHDC15P, VHDC15N, VHDC16P, VHDC16N,
     VHDC17P, VHDC17N, VHDC18P, VHDC18N, VHDC19P, VHDC19N, VHDC20P, VHDC20N
   };
   
// Probes of internal signals:
// Get the FMout signal and clock enables from the VHDC connector:
// These signals are registered internally with the master clock positive edge
wire signed [23:0] FMout       = VHDC[23:0];
wire               clken48kHz  = VHDC[24];
wire               clken192kHz = VHDC[25];
wire               clock_ok    = VHDC[26];

// The data and clock to the external DAC (unsigned data):
wire [6:0] DACdata = {PMOD10, PMOD3, PMOD9, PMOD2, PMOD8, PMOD1, PMOD7};
wire       DACclock = PMOD4;

// Define bit vectors for the buttons, switches and leds:
assign {btnu, btnr, btnd, btnl, btnc} = btns;
assign { sw7, sw6, sw5, sw4, sw3, sw2, sw1, sw0} = sws;
assign leds = { ld7, ld6, ld5, ld4, ld3, ld2, ld1, ld0};

// Local signals for local UART connection:
reg             uart_txen;
wire            uart_rxready, uart_txready;
reg  [7:0]      uart_din;
wire [7:0]      uart_dout;

// Signals to connect to the virtual in/outs of the LM4550 verification IP:
reg  signed [17:0]     LEFT_IN, RIGHT_IN;
wire signed [17:0]     LEFT_OUT, RIGHT_OUT;


//----------------------------------------------------
// UART 921600 baud, 8 bit, 1 stop bit, no parity:
uart   #(
                .INPUT_CLOCK_FREQUENCY( CLOCK_FREQUENCY ), 
                .TX_BAUD_RATE( 921_600 ),
		        .RX_BAUD_RATE( 921_600 )
		)
      uart_sim_1 
	           ( 
				  .clock( BIT_CLK ),	// use the same clock as the codec clock
                  .reset(reset),		// master reset, asynchronous, active high
                  .tx(rx),				// tx data, connected to rx input
                  .rx(tx),				// rx data, connected to tx output
                  .txen(uart_txen),			// load data into transmit buffer and initiate a transmission
                  .txready(uart_txready),	// ready to receive a new byte to tx
                  .rxready(uart_rxready),	// data is ready at dout port
                  .dout(uart_dout),			// data out (received data)
                  .din(uart_din)				// data in (data to transmit)
               );


//----------------------------------------------------
// Simulation model of the LM4550 digital interface:
LM4550_digital_sim  LM4550_digital_sim_1(
            .XTAL_IN( XTAL_IN ),
			.RESET_N( RESET_N ),
			.BIT_CLK( BIT_CLK ),
			.SYNC( SYNC ),
			.SDATA_IN( SDATA_IN ),
			.SDATA_OUT( SDATA_OUT ),
			
			.LEFT_IN( LEFT_IN ),   // inputs to receive the "analogue" audio sent to the ADC
			.RIGHT_IN( RIGHT_IN ), // and transmitted via the AC97 interface
			
			.LEFT_OUT( LEFT_OUT ), // outputs with the "analogue" audio samples from the DAC
			.RIGHT_OUT( RIGHT_OUT )
			);			 
				

//----------------------------------------------------
// Initialize inputs, disable the 100 MHz clock signal (not used in this design):
initial
begin
  // primary inputs:
  clk100M = 1'b0;   // NOT USED !
  btns = 5'b0000_0;
  sws  = 8'b1000_0000;  // Set sw7 to 1 to disable the clock enable generator
  reset_n = 1'b1;
  XTAL_IN = 1'b0;
  
  // to the simulation UART:
  uart_txen = 1'b0;
  uart_din = 8'd0;
end		


// Start the CODEC clock (12.288 MHz). This is the clock source for 
// the system main clock 98.304 MHz
initial
begin
  #2
  forever #( XTAL_PERIOD_NS / 2 ) XTAL_IN = ~XTAL_IN;
end


//------------------------------------------------------
// Generate the external reset signal (note this is active low)
// Activate reset_n for N clock cycles
// The main clock applied to the design is the input clock ( 12.288 MHz )
// multiplied by 8. 
// To avoid racing conditions, reset is delayed 2.6 periods of 98.3 MHz, from the 
// positive edge of XTAL_IN to align the transitions to the negative edge of
// the master internal clock. As we are using a synchronous reset, we must
// wait for the internal clock multiplier to stabilize, otherwise there will be
// no clock to trigger the reset.
//                  ____________________________________________________________________________
// DLL lock _______|
//                    _______________________                         ______________________
//  XTAL_IN  ________|                       |_______________________|                      |__
//(12.288)            __    __    __    __    __    __    __    __    __    __    __    __    _
// 98.3M clk_________|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|
//          __________________________                                                 ________
// reset_n            < --  2.6 T  -->|_______________________..._____________________|
initial
begin
  #1
  // Wait for the DLL lock (clocks running)
  @( posedge clock_ok );
  #1
  @( posedge XTAL_IN );
  # ( 2.6 * INTERNAL_CLOCK_PERIOD );
  reset_n = 1'b0;
  repeat ( N_CLOCKS_RESET )
  begin
    @(negedge XTAL_IN)
    #2;
  end
  reset_n = 1'b1;
end	

// active high reset (used locally only)
assign reset = ~reset_n;


//------------------------------------------------------
// memories for the input and golden output data:
reg signed [17:0]  left_in_mem[ 0: MAX_INPUT_SIZE-1 + 1 ];
reg signed [17:0] right_in_mem[ 0: MAX_INPUT_SIZE-1 + 1 ];

// The output data will be only 24 bit wide
// Samples read from file are 32-bit to simplify the 
// write/read from Matlab and Verilog (???)
reg signed [31:0] FM_golden_out_mem[0:MAX_INPUT_SIZE*4-1 + 1];

// The DAC output golden file:
reg [7:0] DAC_golden_out_mem[0: MAX_INPUT_SIZE*2048-1+1];


// Counts the number of input samples:
integer no_input_samples = 0,
        no_output_samples = 0;

// Counts the number of errors
integer error_count = 0;	

// output file handler:
integer FMfpout, DACfpout;

// Trigger event to start collecting the output data:
event startgetouts;
		
		

//------------------------------------------------------
// Limit the simulation time (maximum number of input samples)
// Use the signal SYNC to count the number of input samples
// coming from the codec
integer clkcount = 0;
always @(posedge SYNC)
begin
  clkcount = clkcount+1;
  if ( clkcount == MAX_SIMULATION_TIME ) 
  begin
    $display("Maximum simulation time exhausted (%d sampling periods).", MAX_SIMULATION_TIME );
	finalize_simulation( );
  end
end


// For plotting in the waveform window:
reg [17:0] error_left=0, error_right=0;

// Set to 1 when the first set of correct samples is detected.
// Verification will only start from that point.
integer start_checking = 0;

// Pointers to vectors:
integer i = 0, j = 0;


//------------------------------------------------------
// Main simulation thread:
initial
begin
  
  // Open text files for output:
  FMfpout  = $fopen( FM_OUTPUT_FILENAME, "w+");  // The FM modultation signal
  DACfpout = $fopen( DAC_OUTPUT_FILENAME, "w+"); // The DAC data

  // Load input datafiles and golden output file:
  $display("Loading simulation input data from files %s, %s:", 
                                     LEFT_IN_FILENAME, RIGHT_IN_FILENAME );
  $readmemh(LEFT_IN_FILENAME,   left_in_mem );
  $readmemh(RIGHT_IN_FILENAME,  right_in_mem );
  
  //-----------------
  // LOAD THE GOLDEN DATA FILES:
  //-----------------
  #1
  // Determine the number of input samples read from files
  // The golden output file will have at least this number of samples x 4:
  no_input_samples = -1;
  for(i=0; i<MAX_INPUT_SIZE; i=i+1)
  begin
    `ifdef DEBUG_PRINT
       if ( i < `NDATA_TO_PRINT )
           $display("Datain(%5d) [ left, right] = [%8d  , %8d] (hex %05H  %05H)", 
		                                                     i, left_in_mem[i], right_in_mem[i],
                                                                left_in_mem[i], right_in_mem[i] );
    `endif
	if ( left_in_mem[i] === 18'dx )
	begin
	  no_input_samples = i;
	  i = MAX_INPUT_SIZE;
	end
  end
  // If read more than MAX_INPUT_SIZE samples...
  if ( no_input_samples == -1 )
    no_input_samples = MAX_INPUT_SIZE;
	
  $display("-----------------------------------------------");
  $display("Read %d samples from input files\n", no_input_samples );
  $display("-----------------------------------------------");
  
  
  
  $display("Loading golden output data from file %s:", FM_GOLDEN_OUTPUT_FILENAME );
  
  // This must be at least 4 X no_input_samples:
  $readmemh( FM_GOLDEN_OUTPUT_FILENAME,  FM_golden_out_mem );
  
  no_output_samples = -1;
  for(i=0; i<MAX_INPUT_SIZE*4; i=i+1)
  begin
    `ifdef DEBUG_PRINT
       if ( i < `NDATA_TO_PRINT )
           $display("Golden dataout(%5d) = %8d (hex %06H )", i, $signed(FM_golden_out_mem[i][23:0]), FM_golden_out_mem[i][23:0] );
    `endif
	if ( FM_golden_out_mem[i] === 32'dx )
	begin
	  no_output_samples = i;
	  i = MAX_INPUT_SIZE*4;
	end
  end
  if ( no_output_samples == -1 )
    no_output_samples = MAX_INPUT_SIZE*4;
	
  $display("-----------------------------------------------");
  $display("Read %d samples from output golden file\n", no_output_samples );
  $display("-----------------------------------------------");
 
  if ( no_output_samples < 4 * no_input_samples )
  begin
    $display("Error: the number of golden samples must be at least equal to 4X the number of input samples");
    $display("Adjusting the number of input samples to %d", no_output_samples/4 );
	no_input_samples = no_output_samples / 4;
    $display("-----------------------------------------------");
  end
  
  // Initialize the "analog" inputs to the CODEC:
  LEFT_IN = 18'd0;
  RIGHT_IN = 18'd0;
    
  # 10
  // wait for the master reset cycle:
  // This will only happen when the master clock is stable:
  @(posedge reset)
  #1
  @(negedge reset);
  #1 
  
  // Program gains of the FM modulator:
  $display("[time=%10.3f us] Reset released, programming gains and output frequency", $time/1000.0 );
  WritePort( { 14'd0, FREQ_STEPWC }  , 8);  // stepWC, freqs 95.50 / 101.60 -> port 8
  WritePort( { 24'd0, GAIN_Kf }, 9);        // Kf = 4     -> port 9
  WritePort( { 28'd0, GAIN_Ks }, 10);       // Ks = 1.000 -> port 10
  WritePort( { 28'd0, GAIN_Kd }, 11);       // Kd = 1.000 -> port 11
  WritePort( { 28'd0, GAIN_Kp }, 12);       // Kp = 0.500 -> port 12
 
  // Wait a few SYNC pulses (input sampling periods) before starting applying the input samples
  // we should receive zeros
  // NOTE: SYNC is generated in the CODEC controller module and is a glitch-free registered output.
  repeat (10)
  begin
	@(posedge SYNC);
	#1;
  end
  
  
  // Start the self-checking verification process:
  -> startgetouts;
  
  
  $display("[time=%10.3f us] Applying input samples...", $time/1000.0 );
  // Apply input samples to the codec "analog" inputs:
  for(i=0; i<no_input_samples; i=i+1 )
  begin
  
    // Start the clock enable generator ONLY when the first data sample arrives to the FM modulator
	if ( i == N_SAMPLES_LATENCY )
	begin
      $display("[time=%10.3f us] Starting the clock enable generator", $time/1000.0 );
      sws[7] = 1'b0; // start clock enable generator
    end
	
    if ( (i % 100 == 0) && (i != 0) )
	  $display("[time=%10.3f us] %5d input samples processed, %3d errors found", $time/1000.0, i, error_count );
	#1
	
	// Apply inputs to the audio CODEC verification model:
    @(posedge SYNC)
	#1;
	LEFT_IN  = left_in_mem[i];
	RIGHT_IN = right_in_mem[i];
	#1;
  end
  
  @(posedge SYNC)
  #1;  
  LEFT_IN  = 18'd0;
  RIGHT_IN = 18'd0; 

  repeat ( 19 )
    @(posedge SYNC)
    
  finalize_simulation( );

end




//------------------------------------------------------
// Self-check process: collect the output of the FM modulator
//  and compare with the golden data:

  // Index to self check golden data vector:
  integer sci = 0;
  
  // Synchronize sampling the output:
  integer synch = 0;
  
  // Loop control variable:
  integer k;
  
  // difference in output and golden values
  integer differror;
  
  // Expected correct data:
  reg [23:0] dataok;
  
  
initial
begin

  // Wait for the event triggered by the input driver:
  @ startgetouts;

  // Discard first output, it will be invalid
  @(negedge clken192kHz );
  #1
  
  // Collect (4 x no_input_samples) output samples:
  for (j=0; j<4*no_input_samples; j=j+1)
  begin
    @(negedge clken192kHz);
	// The FMout output should be directly the output of a register enabled 
	// by the 192 kHz clock enable. 
	// Wait a few clock cycles to probe the output data. As we do not have access to the 
	// master internal clock, we can use the DAC clock to trigger the sampling process:
	repeat (10)
	  @(posedge DACclock);
	
	// Write hex dataout file with the output of the FM modulator:
	$fwrite( FMfpout,"%06h\n", FMout );
	
	// Self check:
	// First we will try to synchronize a match of 5 (?) output samples
	if ( synch == 0 )  // No synch yet, look for the output sample in the first 
	begin              // 5 samples (?) of the golden vector
	  for (k=0; k<10; k=k+1)
	    if ( FMout === FM_golden_out_mem[ k ] && FMout !== 0 ) // Found!
        begin	
		`ifndef DEBUG_PROBES
          $display("Synchronization detected at index %d", k );		
		`endif
		  sci = k;       
		  synch = 1;     // synch found
		  k = 10;        // break loop (tehgere is no 'break' in Verilog ! )
		end
	end
    
    differror = FM_golden_out_mem[ sci ] - FMout ;
	dataok = FM_golden_out_mem[ sci ];
	
	if ( FMout !== FM_golden_out_mem[ sci ] )
	begin
	  `ifdef DEBUG_PRINT
	    `ifndef DEBUG_PROBES
	     if ( j < `NDATA_TO_PRINT*4 )
	     $display("ERROR: Data out (%d) = %d  (%06H), expected %d  (%06H)", j, 
		                                $signed(FMout), $signed(FMout),
										FM_golden_out_mem[ sci ], FM_golden_out_mem[ sci ] );
		 `endif
	  `endif
	  error_count = error_count + 1;
	end
	else
	begin
	  `ifdef DEBUG_PRINT
		 `ifndef DEBUG_PROBES
 	      if ( j < `NDATA_TO_PRINT*4 )
 	        $display("OK:    Data out (%d) = %d  (%06H)", j, $signed(FMout), $signed(FMout) );
		 `endif
	  `endif
	end
	
	sci = sci + 1; // next sample in golden vector
	
  end
  
  finalize_simulation( );
  
end


//------------------------------------------------------
// Virtual register emulates the DAC register:
// Write to hex file:
reg [6:0] DACdataout = 7'd0;
always @(posedge DACclock )
begin
  DACdataout <= DACdata;
  $fwrite( DACfpout,"%02h\n", DACdataout );
end


//------------------------------------------------------
// Check DAC output at each rising clock cycle
initial
begin
  // Wait for the event triggered by the input driver:
  @ startgetouts;

  // Discard first output, it will be invalid
  @(posedge clken192kHz );
  
  while ( 0 )
  begin
    
  end
end


`include "../src/verilog-tb/verilog-tasks.v"

endmodule



