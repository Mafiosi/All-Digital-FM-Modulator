`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:44:22 12/20/2018 
// Design Name: 
// Module Name:    block_sf_192 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module block_sf_192(
	
	input clock,
	input reset,
	input [17:0] LEFT,
	input [17:0] RIGHT,
	output
    );


endmodule
