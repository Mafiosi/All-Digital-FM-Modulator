/*
    Spartan 6 board audio project (V1.4 - Dec 2018)
	
    jca@fe.up.pt

	This Verilog code is property of University of Porto
	Its utilization beyond the scope of the course Digital Systems Design
	(Projeto de Sistemas Digitais) of the Integrated Master in Electrical 
	and Computer Engineering requires explicit authorization from the author.
	
*/

`timescale 1ns/1ps

// Define the module to instantiate:

// Comment next line to instantiate your module:
//`define REFERENCE_MODEL

// Uncomment next line to instantiate your module:
`define  MY_DESIGN    "../src/verilog-rtl/alunos/joaobeleza-pedrocosta/instance.v"


module s6base( 
			//------------------------------------------------------------------
			// Gobal external signals:
			input clockext100MHz,	  // master clock input (external oscillator 100MHz) THIS CLOCK IS NOT USED IN THIS PROJECT
			//------------------------------------------------------------------
			
			input reset_n,            // external reset, active low
			//------------------------------------------------------------------
            // push buttons: button down = logic 1 (no debouncing hw)
			input btnu,			  // button up
			input btnr,           // button right
			input btnd,           // button down
			input btnl,			  // button left
			input btnc,           // button center

			//------------------------------------------------------------------
            // Slide switches:
			input sw0,
			input sw1,
			input sw2,
			input sw3,
			input sw4,
			input sw5,
			input sw6,
			input sw7,

			//------------------------------------------------------------------
			// LEDs: logic 1 lights the LED
			output ld7,			// LED 7 (leftmost)
			output ld6,
			output ld5,
			output ld4,
			output ld3,
			output ld2,
			output ld1,
			output ld0,			// LED 6 (rightmost)


			//------------------------------------------------------------------
			// Serial interface (RS232 port)
            output tx,		// tx data (output from the user circuit)
            input  rx,		// rx data (input to the user circuit)
								
								
			//------------------------------------------------------------------
			// Audio codec interface (LM4550)
			input  SDATA_IN,    // serial stream from codec
			output SDATA_OUT,   // serial stream to codec
			output SYNC,        // frame sync
			input  BIT_CLK,     // bit clock (12.288 MHz)
			output RESET_N,     // codec hw reset (active low)
			
			
			//------------------------------------------------------------------
			// PMOD connector
			output reg PMOD1,  
			output reg PMOD2,  
			output reg PMOD3,  
			output     PMOD4,  
			output reg PMOD7,  
			output reg PMOD8,  
			output reg PMOD9,  
			output reg PMOD10,

			output    VHDC1P,
			output    VHDC1N,
			output    VHDC2P,
			output    VHDC2N,
			output    VHDC3P,
			output    VHDC3N,
			output    VHDC4P,
			output    VHDC4N,
			output    VHDC5P,
			output    VHDC5N,
			output    VHDC6P,
			output    VHDC6N,
			output    VHDC7P,
			output    VHDC7N,
			output    VHDC8P,
			output    VHDC8N,
			output    VHDC9P,
			output    VHDC9N,
			output    VHDC10P,
			output    VHDC10N,
			output    VHDC11P,
			output    VHDC11N,
			output    VHDC12P,
			output    VHDC12N,
			output    VHDC13P,
			output    VHDC13N,
			output    VHDC14P,
			output    VHDC14N,
			output    VHDC15P,
			output    VHDC15N,
			output    VHDC16P,
			output    VHDC16N,
			output    VHDC17P,
			output    VHDC17N,
			output    VHDC18P,
			output    VHDC18N,
			output    VHDC19P,
			output    VHDC19N,
			output    VHDC20P,
			output    VHDC20N
			
			);
								
// VHDC bus (for routing signals to primary outputs):
// assign unused outputs to zero.
wire [39:0] VHDC;
assign 
   { VHDC1P,  VHDC1N, VHDC2P, VHDC2N, VHDC3P, VHDC3N, VHDC4P, VHDC4N, 
     VHDC5P,  VHDC5N, VHDC6P, VHDC6N, VHDC7P, VHDC7N, VHDC8P, VHDC8N, 
     VHDC9P,  VHDC9N,  VHDC10P, VHDC10N, VHDC11P, VHDC11N, VHDC12P, VHDC12N,
     VHDC13P, VHDC13N, VHDC14P, VHDC14N, VHDC15P, VHDC15N, VHDC16P, VHDC16N,
     VHDC17P, VHDC17N, VHDC18P, VHDC18N, VHDC19P, VHDC19N, VHDC20P, VHDC20N
   } = VHDC;

//---------------------------------------------------
// global synchronous reset, active high
reg			reset_d, reset;

//---------------------------------------------------
// UART local signals:
wire        txen, rxready, txready;

//---------------------------------------------------
// data bus between UART and the I/O ports module:
wire [ 7:0] din, dout;

//---------------------------------------------------
// General 32-bit I/O ports:
// output ports (32 bits)
wire [31:0] P0out, P1out, P2out, P3out,
            P4out, P5out, P6out, P7out,
			P8out, P9out, PAout, PBout,
			PCout, PDout, PEout, PFout; 
// input ports (32 bits)			
wire [31:0] P0in,  P1in,  P2in,  P3in,
            P4in,  P5in,  P6in,  P7in;  
				
// Local clocks, generated by the codec, double of the bit clock 12.288 MHz:
// Not used in 2018/2019 project
wire    clock24576k, clock12288k;

// keep reset active while DLL is not locked:
wire clock_ok;


// 
wire clock196M, clock196M_ubf;
wire ckdummy;



// DCM/CMT: receives the 12.288 clock from the CODEC and
// generates the 24.576 and 12.288 main clocks.
// Output "LOCKED" is asserted when the DCM starts generating the 
// clock signal.
clock_bit2x clock_bit2x_1
   (
    .bit_clk_in( BIT_CLK ),          // IN
    // Clock out ports
    .bit_clk_sync( clock12288k ),    // OUT
    .clock24576K( clock24576k ),     // OUT
	 .clock196M( clock196M ), 
	 .ckdummy( ckdummy ),             // unused OUT
    .LOCKED( clock_ok )
	); 	


reg DACclock = 0;
wire clock98MHz;

// Main clock buffer:
BUFG clk98Mbuf( .I( DACclock ), .O( clock98MHz ) );



//---------------------------------------------------
// Reset synchronizer: keep reset active while DDL is not locked:
always @(posedge clock98MHz )
begin
  if ( ~clock_ok )
  begin
    reset <= 1'b1;
  end
  else
  begin
    reset_d <= ~reset_n;
    reset   <= reset_d;
  end
end



//---------------------------------------------------
// UART 921600 baud, 8 bit, 1 stop bit, no parity:
uart  #( 
         .INPUT_CLOCK_FREQUENCY( 98_304_000 ),
         .TX_BAUD_RATE( 921_600 ),
		   .RX_BAUD_RATE( 921_600 )
		)
        uart_1 
 		   ( 
             .clock( clock98MHz ),	// master clock (100MHz)
             .reset(reset),			// master reset, asynchronous, active high
             .tx(tx),					// tx data, connected to rx input
             .rx(rx),					// rx data, connected to tx output
             .txen(txen),			// load data into transmit buffer and initiate a transmission
             .txready(txready),	// ready to receive a new byte to tx
             .rxready(rxready),	// data is ready at dout port
             .dout(dout),			// data out (received data)
             .din(din)				// data in (data to transmit)
           );

//---------------------------------------------------
// Command interpreter:
ioports16V2018
            #(   // Define initial reset values for the output ports (default is 32'd0)
                 .INIT_P08( { 14'd0, 18'b000010001001010100 } ), // Stepwc = 2.145263671875 (FM freqs  95.00 MHz and 101.60 MHz)
                 .INIT_P09( { 24'd0,  8'b0100_0000 } ),			 // Kf = 4.000
                 .INIT_P10( { 28'd0,  4'b1000 } ),               // Ks = 1.000
                 .INIT_P11( { 28'd0,  4'b1000 } ),			     // Kd = 1.000
                 .INIT_P12( { 28'd0,  4'b0100 } ) 	             // Kp = 0.500
             )

// ioports
 				 ioports16_1 
             ( 
			      .clk( clock98MHz ),	// master clock 
               .reset(reset),		   // master reset, asynchronous, active high
               
               .load(rxready),		// load enable for din bus
               .ready(txready),		// ready to consume dout data
               .enout(txen),		   // enable loading of dout data
               
               .datain(dout),		// data in bus (8 bits), from USART
               .dataout(din),		// data out bus (8 bits), to USART
               
               .in0(P0in),	.in1(P1in), .in2(P2in), .in3(P3in),
					.in4(P4in), .in5(P5in), .in6(P6in), .in7(P7in),			
               
               .out0(P0out), .out1(P1out), .out2(P2out), .out3(P3out),			 
			      .out4(P4out), .out5(P5out), .out6(P6out), .out7(P7out),
			      .out8(P8out), .out9(P9out), .outa(PAout), .outb(PBout),
			      .outc(PCout), .outd(PDout), .oute(PEout), .outf(PFout)
			);
					
					
//---------------------------------------------------------------------------------
// LM5440 audio CODEC interface
wire [15:0]DIN;
wire [5:0] REGID;
wire [3:0] STATUS;
wire WE, RE, RDY, DIN_RDY, DOUT_RQST;

wire [17:0] LEFT_in, RIGHT_in,      // From the codec
            LEFT_inf, RIGHT_inf,    // After selector controlled by sw5/sw4 to ground left or right channels
            LEFT_out, RIGHT_out;    // To codec; sw7/sw6 select to the codec the outputs from the filters of the inputs			

LM4550_controler LM4550_controler_1 (
                .SDATA_IN(SDATA_IN),
                .SDATA_OUT(SDATA_OUT),
                .SYNC(SYNC),
                .BIT_CLK( clock12288k ),        // bit clock 12.288 MHz
                .RESET_N( ),                    // Reset to external codec
                .DIN(DIN),
                .REGID(REGID),
                .STATUS(STATUS),
                .WE(WE),
                .RE(RE),
                .RDY(RDY),
					 
                .DIN_RDY(DIN_RDY),          // Data input enable
                .RIGHT_IN( RIGHT_in ),      // from codec
                .LEFT_IN( LEFT_in ),
					 
                .DOUT_RQST(DOUT_RQST),     // request for output data to DAC
                .RIGHT_OUT( RIGHT_out ),   // to codec
                .LEFT_OUT( LEFT_out ),
					 
                .RESET(reset),
                .CLOCK( clock98MHz )
				);
				
// Disable CODEC reset:				
assign RESET_N = 1'b1;				
					 
// assign control signals to access the LM4550 programming interface:					 
assign DIN=P2out[15:0];
assign REGID=P3out[5:0];
assign P1in={27'b0,STATUS};
assign WE=PFout[0];
assign RE=PFout[1];
assign P2in={31'd0,RDY};


// Synchronize the audio data coming from the CODEC to the local 48k clock enable

// Delay the DIN_RDY signal by 3 clock cycles:
reg [2:0] r_dinrdy;
always @(posedge clock98MHz )
if ( reset )
begin
  r_dinrdy <= 3'b000;
end
else
begin
  r_dinrdy <= { r_dinrdy[1:0], DIN_RDY };
end

// This is the                                                                                                                                                                                                                                         clock enable 48 kHz generated by the audio codec controller:
wire   din_en;
assign din_en = ~r_dinrdy[1] & r_dinrdy[2];


// Clock enable generator. This is required to guarantee the 
// relative timing between the two clock enable signals
wire clken48kHz_c, clken192kHz_c;
reg  clken48kHz,   clken192kHz;
wire run_genclock;
assign run_genclock = ~sw7;
clockenablegen clken48k192k( 
                .clock( clock98MHz ),
			    .reset( reset ),
				.run( run_genclock ),
			    .clken48kHz( clken48kHz_c ),
			    .clken192kHz( clken192kHz_c )
			);
					 
					 
// Audio databus synchronized to the user 48 kHz clock enable:
reg signed [17:0] leftins, rightins;
always @(posedge clock98MHz )
if ( reset )
begin
  leftins  <= 18'd0;
  rightins <= 18'd0;
  clken48kHz <= 1'b0;
  clken192kHz <= 1'b0;
end
else
begin
  if ( clken48kHz_c )
  begin
    leftins  <= LEFT_in;
    rightins <= RIGHT_in;
  end
  clken48kHz <= clken48kHz_c;
  clken192kHz <= clken192kHz_c;
end

					 
//-------------------------------------------------------------------------------
// Audio samples are available in the positive clock edge when din_en is 1
// 
// A synchronous process to handle the audio stream should be as:
// always @(posedge clock)
// if ( reset )
//   // do the reset actions
// else
//   if ( din_en )
//   begin
//     // do something with rightins and leftins
//     // and generate rightouts and leftouts
//   end
//-------------------------------------------------------------------------------


//-------------------------------------------------------------------------------
// Implement some basic functions using  the audio stream
// The modulation signal (see below)
reg signed [13:0] datamod;
//
// Set sw0=1 / sw1=1  to mute left/right inputs:
// set sw2=1 / sw3=1 to swap left and right channels
assign LEFT_inf   = ( sw0 ) ? 18'd0 : ( sw2 ? rightins : leftins  );
assign RIGHT_inf  = ( sw1 ) ? 18'd0 : ( sw3 ? leftins  : rightins );	

assign LEFT_out   = LEFT_in;					 
assign RIGHT_out  = RIGHT_in;	
			 				 				 
// Generate the output mono signal rectified to view the mono signal envelope:
wire [18:0] mono_digital_mix;
wire [18:0] mono_digital_mix_rectified;
assign mono_digital_mix =  ( {LEFT_inf[17], LEFT_inf} + {RIGHT_inf[17], RIGHT_inf} ) / 2;
assign mono_digital_mix_rectified = mono_digital_mix[17] ? ( -mono_digital_mix ) : ( mono_digital_mix );	


//-------------------------------------------------------------------------------
// display the output signal envelope
assign {ld7, ld6, ld5, ld4, ld3, ld2, ld1, ld0} = mono_digital_mix_rectified[18:11];  
  

//-------------------------------------------------------------------------------
// Generate the DAC clock using the double frequency clock (2 x 98.304 MHz)
always  @( posedge clock196M )
begin
  DACclock <= ~DACclock;
end

//-------------------------------------------------------------------------------  
// Connect the DAC clock to the PMOD output (connector pin 4)
assign PMOD4 = DACclock;


//-------------------------------------------------------------------------------  
// Connect the datapath gains:
wire        [7:0] Kf;
wire        [3:0] Ks, Kd, Kp;
assign Kf = P9out[7:0];  // Port 9
assign Ks = PAout[3:0];  // Port 10
assign Kd = PBout[3:0];  // Port 11
assign Kp = PCout[3:0];  // Port 12

wire signed [23:0] FMout;


`ifdef REFERENCE_MODEL
//-------------------------------------------------------------------------------  
// Instgantiate the FM stereo modulator
stereo_fm_mx_golden  stereo_fm_mx_golden_1(
				//-----------------------------------------------
				// Global signals
                .clock( clock98MHz ),     // master clock, active in posedge
                .reset( reset ),     // master reset, synchronous, active high
				
				//-----------------------------------------------
				// Gains:
				.Ks( Ks ),
				.Kd( Kd ),
				.Kp( Kp ),
				.Kf( Kf ),
				//-----------------------------------------------
			
				//-----------------------------------------------
				// Audio data in:
               .LEFTin( LEFT_inf ),            // data in, left channel
               .RIGHTin( RIGHT_inf ),          // data in, right channel

				.clken48kHz( clken48kHz ),    // Clock enable for input sampling rate:
				.clken192kHz( clken192kHz ),  // Clock enable for 4X sampling rate:
				
				//-----------------------------------------------
				// FM Stereo dataout:
				.FMout( FMout )               // data out, FM stereo signal
            );


`endif

`ifdef MY_DESIGN
  `include `MY_DESIGN
`endif


//-------------------------------------------------------------------------------  
// Generate the modulation signal
// Test signal to modulate: 14 bits, signed:

//-------------------------------------------------------------------------------  
// Generate a test signal (central "LA" = 440 Hz)
wire signed [7:0] test440Hz;
//ddsaudio #( .OUTPUT_FREQUENCY( 440 ) 
//          )
ddsaudio		  dds_test_signal
		  (
		.clock( clock98MHz ),
		.reset( reset ),
		.enableclk( clken48kHz ),
		.outsine( test440Hz )
        );


reg signed [13:0] testmod; 
reg signed [15:0] testmodlong;


always @(posedge clock98MHz )
begin
  if ( reset )
  begin
    testmodlong  <= 0;
    testmod      <= 0;
    datamod      <= 0;
  end
  else
  begin
	// testmod = 8 bit sine wave + 8 bit gain kf = 16 bits >> 2 = 14 bits
    testmodlong  <= ( $signed( test440Hz ) * $signed( { 1'b0, Kf }) ); 
    testmod      <= testmodlong >>> 2;
	 
    datamod      <= sw6 ? testmod : FMout[23:10];  
  end
end


//-------------------------------------------------------------------------------  
// output the FMout signal and clock enables to the VHDC connector:
reg [23:0] FMout_r;
reg        clken48kHz_r;
reg        clken192kHz_r;

always @(posedge clock98MHz )
begin
  if ( reset )
  begin
    FMout_r        <= 0;
    clken48kHz_r   <= 0;
    clken192kHz_r  <= 0;
  end
  else
  begin
    FMout_r        <= FMout      ;
    clken48kHz_r   <= clken48kHz ;
    clken192kHz_r  <= clken192kHz;
  end
end

assign VHDC[23:0] = FMout_r;
assign VHDC[24]   = clken48kHz;
assign VHDC[25]   = clken192kHz;
assign VHDC[26]   = clock_ok;
// connect to zero the unused VHDC outputs:
assign VHDC[39:27] = 0;


//-------------------------------------------------------------------------------  
// Connect the phase step input to tune the output frequency:
wire signed [19:0] stepwc;
assign stepwc = P8out[19:0];


//-------------------------------------------------------------------------------  
// The final DDS
wire [7:0] datasine;
dds_carrier dds_carrier_1(
        .clock( clock98MHz ),
        .reset( reset ),
		.enableclk( 1'b1 ),
		.phasein( datamod ),
		.stepwc( stepwc ),
		.outsine( datasine )
    );


// Data to the external DAC:
reg [6:0] dataDAC;
always  @( posedge clock98MHz )
if ( reset ) 
begin
  dataDAC <= 7'b0;
end
else
begin
  // datasine is signed but the DAC requires unsigned data:
  dataDAC <= { ~datasine[7], datasine[6:1] };
end


//--------------------------------------------------
// Connect to the DAC inputs:
// PMOD connector (front view)
//  Vcc  GND    CLK  D8   D6   D4
//   6    5      4    3    2    1 <<-- PMOD pin number
//   O    O      O    O    O    O
//   O    O      O    O    O    O
//  12   11     10    9    8    7 <<-- PMOD pin number
//  Vcc  GND    D9   D7   D5   D3
//

always @ (posedge clock98MHz ) // 98 MHz
if ( reset )
begin
  {PMOD10, PMOD3, PMOD9, PMOD2, PMOD8, PMOD1, PMOD7} <= 7'd0;
end
else
begin
  {PMOD10, PMOD3, PMOD9, PMOD2, PMOD8, PMOD1, PMOD7} <= dataDAC;
end


  


//---------------------------------------------------------------------------------
// Connect P0in to the push buttons and slide switches:
assign P0in[31:21] = 32'd0;
assign P0in[20:16] = {btnu, btnr, btnd, btnl, btnc };
assign P0in[15: 8] = 8'd0;
assign P0in[ 7: 0] = {sw7, sw6, sw5, sw4, sw3, sw2, sw1, sw0};

// Unused input ports
assign P3in[31:24]  = 32'd0;
assign P4in[31:18]  = 32'd0;
assign P5in[31:24]  = 32'd0;
assign P6in[31:24]  = 32'd0;
assign P7in[31:24]  = 32'd0;
//---------------------------------------------------------------------------------


		
endmodule

