//-------------------------------------------------------------------------------
//  FEUP / MIEEC - Digital Systems Design 2018/2019
//
//  Module for Lab Project 3: 
//     Implementation of an All-digital FM stereo Modulator
//  
//  MIEEC - Jo�o Beleza up201402831@fe.up.pt
//          Pedro Costa up201402793@fe.up.pt
//
//  DELIVER DATE: XX/XX/201X
//-------------------------------------------------------------------------------

`timescale 1ns / 1ps

module Lin_inter(
	 input clock,
	 input reset,
    input [17:0] LI_mR_in,
    input [17:0] LI_pR_in,
    output [17:0] LI_mR_out,
    output [17:0] LI_pR_out
    );


endmodule
